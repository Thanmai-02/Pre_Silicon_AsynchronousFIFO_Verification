typedef uvm_sequencer#(read_transaction) read_sequencer;