typedef uvm_sequencer#(write_transaction) write_sequencer;